module alu_mov(
  input wire  [15:0] operand1,
  output wire  [15:0] dout);
  
  assign dout = operand1;
  
endmodule 